Star Wars är en franchise som främst består av en serie amerikanska science fiction-filmer skapade av George Lucas under 1970-, 1980-, 1990-, 2000- och 2010-talet. Den första i filmserien, Stjärnornas krig, hade premiär 25 maj 1977 i 
USA och blev snabbt ett världsomfattande populärkulturfenomen. Filmens framgång ledde till två uppföljare, Rymdimperiet slår tillbaka (1980) och Jedins återkomst (1983). Tjugotvå år efter den ursprungliga filmens premiär började George 
Lucas arbetet med en andra trilogi som en prequel till originaltrilogin bestående av Episod I – Det mörka hotet (1999), Episod II – Klonerna anfaller (2002) och Episod III – Mörkrets hämnd (2005). Under 2012 sålde Lucas 
rättigheterna till Walt Disney Company. Tio år efter Episod III släpptes den första delen i uppföljartrilogin, den sjunde filmen i serien Episod VII – The Force Awakens (2015). Ytterligare två uppföljare är planerade, Episod VIII 
(2017) och Episod IX (2019).

Filmserien har också resulterat i böcker, tv-serier, datorspel och serietidningar. Dessa tillägg utgör grunden för Star Wars: Expanded Universe, och har resulterat i en märkbar utveckling i seriens fiktiva universum. Fram till mars 
2016 har de sex filmerna tillsammans genererat uppskattningsvis 9,2 miljarder US dollar, vilket gör dem till den tredje mest inkomstbringande filmserien.[1]
